`timescale 1ns / 1ps
/*
 * The MIT License (MIT)
 *
 * Copyright (c) 2015 Robert Armstrong
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 * 
 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

module mdio_1to2
    (input  wire mdio_mdc,
     input  wire mdio_o,
     input  wire mdio_t,
     output wire mdio_i,

     output wire phy0_mdc,
     output wire phy0_mdio_o,
     output wire phy0_mdio_t,
     input  wire phy0_mdio_i,

     output wire phy1_mdc,
     output wire phy1_mdio_o,
     output wire phy1_mdio_t,
     input  wire phy1_mdio_i
     );

    assign phy0_mdc    = mdio_mdc;
    assign phy0_mdio_t = mdio_t;
    assign phy0_mdio_o = mdio_o;

    assign phy1_mdc    = mdio_mdc;
    assign phy1_mdio_t = mdio_t;
    assign phy1_mdio_o = mdio_o;

    assign mdio_i      = phy0_mdio_i & phy1_mdio_i;

endmodule
